package Hard_Update2.0_pkg;

// =============================================================================
// Generated Register Block 1.0
// Commit ID: aa9d7e6ebfe1c3a5f842cb190dfae6cd73d7e4fa
// =============================================================================

typedef struct packed {
  logic [31: 0] wptr;
} WPTR_t;

typedef struct packed {
  logic [31: 0] fetch_rptr;
} FETCH_RPTR_t;

endpackage : Hard_Update2.0_pkg
