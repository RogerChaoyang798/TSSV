package AIGC_DEMO_reg_pkg;

// =============================================================================
// Register bit field definition
// =============================================================================

