import Hard_Update2.0_pkg::*;

// =============================================================================
// Generated Register Block 1.0
// =============================================================================

                
               
        module Hard_Update2.0 
           (
           input   clk,
   input   rst_b,
   input  [11:0] paddr,
   input  [31:0] pwdata,
   output  [31:0] prdata,
   input   psel,
   input   penable,
   input   pwrite,
   output   pready,
   output reg   pslverr,
   output  [31:0] cfg_wptr,
   input   wptr_update,
   input  [31:0] wptr_update_value,
   output  [31:0] cfg_fetch_rptr,
   input   fetch_rptr_update,
   input  [31:0] fetch_rptr_update_value
           );
        
           wire  reg_rd;
   wire  reg_wr;
   wire [11:0] reg_addr;
   reg [31:0] reg_rdata;
   wire [31:0] reg_wdata;
   wire [31:0] next_rdata;
   wire  in_range;
   wire  slverr;
   wire  dec_wptr;
   reg [31:0] reg_wptr;
   wire  wptr_we;
   wire  dec_fetch_rptr;
   reg [31:0] reg_fetch_rptr;
   wire  fetch_rptr_we;
        
        // apb interface
assign prdata = reg_rdata;
assign reg_wr = psel && penable && pwrite;
assign reg_rd = psel && !penable && !pwrite;
assign pready = 1'b1;
assign slverr = psel && !in_range;
assign reg_addr = paddr;
assign reg_wdata = pwdata;
assign dec_wptr = (reg_addr == 12'hF000) ? 1'd1 : 1'd0;
assign wptr_we = reg_wr && dec_wptr;
// non-RO: output
assign cfg_wptr = reg_wptr;
assign dec_fetch_rptr = (reg_addr == 12'hF004) ? 1'd1 : 1'd0;
assign fetch_rptr_we = reg_wr && dec_fetch_rptr;
// non-RO: output
assign cfg_fetch_rptr = reg_fetch_rptr;
assign in_range = |{dec_wptr,
dec_fetch_rptr};
// Read data mux
assign next_rdata = 
( {32{dec_wptr}} & reg_wptr ) |
( {32{dec_fetch_rptr}} & reg_fetch_rptr );

    
        
    
        
always @( posedge clk  or negedge rst_b )

       if(!rst_b)
       begin
    pslverr <= 1'h0;
      end
  else
  begin
  pslverr <= slverr;
  end
  

always @( posedge clk  or negedge rst_b )

       if(!rst_b)
       begin
    reg_wptr <= 32'h0;
      end
  else if(wptr_we)
  begin
  reg_wptr <= reg_wdata;
  end
  else if(wptr_update)
  begin
  reg_wptr <= wptr_update_value;
  end
  

always @( posedge clk  or negedge rst_b )

       if(!rst_b)
       begin
    reg_fetch_rptr <= 32'h0;
      end
  else if(fetch_rptr_we)
  begin
  reg_fetch_rptr <= reg_wdata;
  end
  else if(fetch_rptr_update)
  begin
  reg_fetch_rptr <= fetch_rptr_update_value;
  end
  

always @( posedge clk  or negedge rst_b )

       if(!rst_b)
       begin
    reg_rdata <= 32'h0;
      end
  else if(reg_rd)
  begin
  reg_rdata <= next_rdata;
  end
  

        
        endmodule
         : Hard_Update2.0
